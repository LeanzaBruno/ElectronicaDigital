library ieee;
use ieee.std_logic_1164.all;


entity codificador_tb is
  port
